`ifndef FrameCoprocessor_v1_0_tb_include_vh_
`define FrameCoprocessor_v1_0_tb_include_vh_

//Configuration current bd names
`define BD_NAME FrameCoprocessor_v1_0_bfm_1
`define BD_INST_NAME FrameCoprocessor_v1_0_bfm_1_i
`define BD_WRAPPER FrameCoprocessor_v1_0_bfm_1_wrapper

//Configuration address parameters
`endif
